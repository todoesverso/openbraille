* EESchema Netlist Version 1.1 (Spice format) creation date: 13/1/2009-21:00:19


U1  30 0 2 7805
C1  30 0 0.1u
C2  2 0 0.1u
R6  23 2 3k3
D1  23 0 LED
C4  24 0 10u
U***1  7 18 28 3 0 15 16 14 27 25 26 24 19 2 4 29 22 11 PIC16F84A
X1  29 4 4MHz
RV1  5 2 2 POT10k
C5  0 4 33p
C6  29 0 33p
R4  3 2 10k
SW2  0 3 RESET
Q3  0 17 21 TIP122
K1  2 0 30 CONN_3
R5  5 24 1k
R11  6 22 3k3
R10  12 11 3k3
R9  17 7 3k3
R8  13 18 3k3
SW1  15 0 Left
SW3  14 0 Right
SW4  16 0 Stop
R3  14 2 10k
R2  16 2 10k
R1  15 2 10k
R7  10 19 3k3
Q1  0 10 24 BC337
P1  30 9 21 8 20 0 CONN_6
Q2  0 13 9 TIP122
Q4  0 12 8 TIP122
Q5  0 6 20 TIP122
C3  30 0 100u

.end
